import uvm_pkg::*;

`include "uvm_macros.svh"

`include "dut/apb_if.sv"


`include "testbench/transaction.sv"
`include "testbench/reg.sv"
`include "testbench/reg_block.sv"
`include "testbench/adapter.sv"
`include "testbench/driver.sv"
`include "testbench/monitor.sv"
`include "testbench/agent.sv"
`include "testbench/scoreboard.sv"
`include "testbench/env.sv"
`include "testbench/reg_sequence.sv"
`include "testbench/test.sv"


`include "dut/apb.sv"